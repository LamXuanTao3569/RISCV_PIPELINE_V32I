module decode_cycle(clk, rst, InstrD, PCD, PCPlus4D, RegWriteW, RDW, ResultW, RegWriteE, ALUSrcE, MemWriteE, ResultSrcE, StallD, FlushD, Jump,
    BranchE,  ALUControlE, RD1_E, RD2_E, Imm_Ext_E, RD_E, PCE, PCPlus4E, RS1_E, RS2_E);

    // Declaring I/O
    input clk, rst, RegWriteW, StallD, FlushD; // Thêm StallD, FlushD
    input [4:0] RDW;
    input [31:0] InstrD, PCD, PCPlus4D, ResultW;

    output RegWriteE,ALUSrcE,MemWriteE,BranchE,Jump;
	 output [1:0] ResultSrcE; // Mở rộng thành [1:0]
    output [2:0] ALUControlE;
    output [31:0] RD1_E, RD2_E, Imm_Ext_E;
    output [4:0] RS1_E, RS2_E, RD_E;
    output [31:0] PCE, PCPlus4E;

    // Declare Interim Wires
    wire RegWriteD, ALUSrcD, MemWriteD, BranchD, JumpD; // Thêm JumpD
    wire [1:0] ResultSrcD; // Mở rộng thành [1:0]
    wire [2:0] ImmSrcD; // Mở rộng thành [2:0]
    wire [2:0] ALUControlD;
    wire [31:0] RD1_D, RD2_D, Imm_Ext_D;

    // Declaration of Interim Register
    reg RegWriteD_r, ALUSrcD_r, MemWriteD_r, BranchD_r, JumpD_r; // Thêm JumpD_r
    reg [1:0] ResultSrcD_r; // Mở rộng thành [1:0]
    reg [2:0] ALUControlD_r;
    reg [31:0] RD1_D_r, RD2_D_r, Imm_Ext_D_r;
    reg [4:0] RD_D_r, RS1_D_r, RS2_D_r;
    reg [31:0] PCD_r, PCPlus4D_r;


    // Initiate the modules
    // Control Unit
    Control_Unit_Top control (
                            .Op(InstrD[6:0]),
                            .RegWrite(RegWriteD),
                            .ImmSrc(ImmSrcD),
                            .ALUSrc(ALUSrcD),
                            .MemWrite(MemWriteD),
                            .ResultSrc(ResultSrcD),
                            .Branch(BranchD),
									 .Jump(JumpD), // Thêm JumpD
                            .funct3(InstrD[14:12]),
                            .funct7(InstrD[31:25]),
                            .ALUControl(ALUControlD)
                            );

    // Register File
    Register_File rf (
                        .clk(clk),
                        .rst(rst),
                        .WE3(RegWriteW),
                        .WD3(ResultW),
                        .A1(InstrD[19:15]),
                        .A2(InstrD[24:20]),
                        .A3(RDW),
                        .RD1(RD1_D),
                        .RD2(RD2_D)
                        );

    // Sign Extension
    Sign_Extend extension (
                        .In(InstrD[31:0]),
                        .Imm_Ext(Imm_Ext_D),
                        .ImmSrc(ImmSrcD)
                        );

    // Declaring Register Logic
    always @(posedge clk or negedge rst) begin
        if(rst == 1'b0) begin
            RegWriteD_r <= 1'b0;
            ALUSrcD_r <= 1'b0;
            MemWriteD_r <= 1'b0;
            ResultSrcD_r <= 1'b0;
            BranchD_r <= 1'b0;
				JumpD_r <= 1'b0; // Thêm JumpD_r
            ALUControlD_r <= 3'b000;
            RD1_D_r <= 32'h00000000; 
            RD2_D_r <= 32'h00000000; 
            Imm_Ext_D_r <= 32'h00000000;
            RD_D_r <= 5'h00;
            PCD_r <= 32'h00000000; 
            PCPlus4D_r <= 32'h00000000;
            RS1_D_r <= 5'h00;
            RS2_D_r <= 5'h00;
        end
		  else if (StallD) begin // Thêm StallD
            // Giữ nguyên giá trị nếu stall
        end
        else begin
            RegWriteD_r <= FlushD ? 1'b0 : RegWriteD;
            ALUSrcD_r <= FlushD ? 1'b0 : ALUSrcD;
            MemWriteD_r <= FlushD ? 1'b0 : MemWriteD;
            ResultSrcD_r <= FlushD ? 2'b00 : ResultSrcD;
            BranchD_r <= FlushD ? 1'b0 : BranchD;
            JumpD_r <= FlushD ? 1'b0 : JumpD;
            ALUControlD_r <= FlushD ? 3'b000 : ALUControlD;
            RD1_D_r <= FlushD ? 32'h00000000 : RD1_D; 
            RD2_D_r <= FlushD ? 32'h00000000 : RD2_D; 
            Imm_Ext_D_r <= FlushD ? 32'h00000000 : Imm_Ext_D;
            RD_D_r <= FlushD ? 5'h00 : InstrD[11:7];
            PCD_r <= FlushD ? 32'h00000000 : PCD; 
            PCPlus4D_r <= FlushD ? 32'h00000000 : PCPlus4D;
            RS1_D_r <= FlushD ? 5'h00 : InstrD[19:15];
            RS2_D_r <= FlushD ? 5'h00 : InstrD[24:20];
        end
    end

    // Output asssign statements
    assign RegWriteE = RegWriteD_r;
    assign ALUSrcE = ALUSrcD_r;
    assign MemWriteE = MemWriteD_r;
    assign ResultSrcE = ResultSrcD_r;
    assign BranchE = BranchD_r;
	 assign JumpE = JumpD_r; // Thêm JumpE
    assign ALUControlE = ALUControlD_r;
    assign RD1_E = RD1_D_r;
    assign RD2_E = RD2_D_r;
    assign Imm_Ext_E = Imm_Ext_D_r;
    assign RD_E = RD_D_r;
    assign PCE = PCD_r;
    assign PCPlus4E = PCPlus4D_r;
    assign RS1_E = RS1_D_r;
    assign RS2_E = RS2_D_r;

endmodule
