module wb_stage (
    input clk, reset, stall,
    input [31:0] mem_wb_result_in,
    input [4:0] mem_wb_rd_in,
    input mem_wb_reg_write_in
);
    // Không có logic hoặc output thêm
endmodule